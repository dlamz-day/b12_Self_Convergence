module spice_pwr_supply 
(
    //======input======
    
    //======output======
    output vdd,
    output vss
);



endmodule  