##
## LEF for PtnCells ;
## created by Encounter v14.28-s033_1 on Thu Sep 15 16:35:22 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO BISG_TOP
  CLASS BLOCK ;
  SIZE 157.2500 BY 153.7200 ;
  FOREIGN BISG_TOP 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 -0.0700 157.2500 0.0700 ;
    END
  END clk
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 4.5900 157.2500 4.7300 ;
    END
  END rst_n
  PIN k[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 23.2200 157.2500 23.3600 ;
    END
  END k[3]
  PIN k[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 18.5600 157.2500 18.7000 ;
    END
  END k[2]
  PIN k[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 13.9050 157.2500 14.0450 ;
    END
  END k[1]
  PIN k[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 9.2450 157.2500 9.3850 ;
    END
  END k[0]
  PIN nl[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 41.8500 157.2500 41.9900 ;
    END
  END nl[3]
  PIN nl[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 37.1950 157.2500 37.3350 ;
    END
  END nl[2]
  PIN nl[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 32.5350 157.2500 32.6750 ;
    END
  END nl[1]
  PIN nl[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 27.8800 157.2500 28.0200 ;
    END
  END nl[0]
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 46.5100 157.2500 46.6500 ;
    END
  END start
  PIN nloss
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 51.1700 157.2500 51.3100 ;
    END
  END nloss
  PIN speaker
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 55.8250 157.2500 55.9650 ;
    END
  END speaker
  PIN ScanNum[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.1750 0.0000 157.3150 0.5000 ;
    END
  END ScanNum[19]
  PIN ScanNum[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 148.9000 0.0000 149.0400 0.5000 ;
    END
  END ScanNum[18]
  PIN ScanNum[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 140.6200 0.0000 140.7600 0.5000 ;
    END
  END ScanNum[17]
  PIN ScanNum[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 132.3450 0.0000 132.4850 0.5000 ;
    END
  END ScanNum[16]
  PIN ScanNum[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 124.0700 0.0000 124.2100 0.5000 ;
    END
  END ScanNum[15]
  PIN ScanNum[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.7950 0.0000 115.9350 0.5000 ;
    END
  END ScanNum[14]
  PIN ScanNum[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.5200 0.0000 107.6600 0.5000 ;
    END
  END ScanNum[13]
  PIN ScanNum[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.2400 0.0000 99.3800 0.5000 ;
    END
  END ScanNum[12]
  PIN ScanNum[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.9650 0.0000 91.1050 0.5000 ;
    END
  END ScanNum[11]
  PIN ScanNum[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.6900 0.0000 82.8300 0.5000 ;
    END
  END ScanNum[10]
  PIN ScanNum[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.4150 0.0000 74.5550 0.5000 ;
    END
  END ScanNum[9]
  PIN ScanNum[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.1400 0.0000 66.2800 0.5000 ;
    END
  END ScanNum[8]
  PIN ScanNum[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 57.8600 0.0000 58.0000 0.5000 ;
    END
  END ScanNum[7]
  PIN ScanNum[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 49.5850 0.0000 49.7250 0.5000 ;
    END
  END ScanNum[6]
  PIN ScanNum[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 41.3100 0.0000 41.4500 0.5000 ;
    END
  END ScanNum[5]
  PIN ScanNum[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.0350 0.0000 33.1750 0.5000 ;
    END
  END ScanNum[4]
  PIN ScanNum[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.7600 0.0000 24.9000 0.5000 ;
    END
  END ScanNum[3]
  PIN ScanNum[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.4800 0.0000 16.6200 0.5000 ;
    END
  END ScanNum[2]
  PIN ScanNum[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 8.2050 0.0000 8.3450 0.5000 ;
    END
  END ScanNum[1]
  PIN ScanNum[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.0700 0.0000 0.0700 0.5000 ;
    END
  END ScanNum[0]
  PIN ADPLL_LOCK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT -0.0700 153.2200 0.0700 153.7200 ;
    END
  END ADPLL_LOCK
  PIN t_p_dec[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 89.7850 153.2200 89.9250 153.7200 ;
    END
  END t_p_dec[7]
  PIN t_p_dec[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 78.5550 153.2200 78.6950 153.7200 ;
    END
  END t_p_dec[6]
  PIN t_p_dec[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.3200 153.2200 67.4600 153.7200 ;
    END
  END t_p_dec[5]
  PIN t_p_dec[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.0900 153.2200 56.2300 153.7200 ;
    END
  END t_p_dec[4]
  PIN t_p_dec[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 44.8600 153.2200 45.0000 153.7200 ;
    END
  END t_p_dec[3]
  PIN t_p_dec[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 33.6250 153.2200 33.7650 153.7200 ;
    END
  END t_p_dec[2]
  PIN t_p_dec[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 22.3950 153.2200 22.5350 153.7200 ;
    END
  END t_p_dec[1]
  PIN t_p_dec[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 11.1600 153.2200 11.3000 153.7200 ;
    END
  END t_p_dec[0]
  PIN range[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.1800 153.2200 157.3200 153.7200 ;
    END
  END range[5]
  PIN range[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 145.9450 153.2200 146.0850 153.7200 ;
    END
  END range[4]
  PIN range[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.7150 153.2200 134.8550 153.7200 ;
    END
  END range[3]
  PIN range[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.4800 153.2200 123.6200 153.7200 ;
    END
  END range[2]
  PIN range[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.2500 153.2200 112.3900 153.7200 ;
    END
  END range[1]
  PIN range[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.0200 153.2200 101.1600 153.7200 ;
    END
  END range[0]
  PIN pass
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 60.4850 157.2500 60.6250 ;
    END
  END pass
  PIN sig[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 121.0400 157.2500 121.1800 ;
    END
  END sig[12]
  PIN sig[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 116.3800 157.2500 116.5200 ;
    END
  END sig[11]
  PIN sig[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 111.7200 157.2500 111.8600 ;
    END
  END sig[10]
  PIN sig[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 107.0650 157.2500 107.2050 ;
    END
  END sig[9]
  PIN sig[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 102.4050 157.2500 102.5450 ;
    END
  END sig[8]
  PIN sig[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 97.7500 157.2500 97.8900 ;
    END
  END sig[7]
  PIN sig[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 93.0900 157.2500 93.2300 ;
    END
  END sig[6]
  PIN sig[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 88.4300 157.2500 88.5700 ;
    END
  END sig[5]
  PIN sig[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 83.7750 157.2500 83.9150 ;
    END
  END sig[4]
  PIN sig[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 79.1150 157.2500 79.2550 ;
    END
  END sig[3]
  PIN sig[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 74.4600 157.2500 74.6000 ;
    END
  END sig[2]
  PIN sig[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 69.8000 157.2500 69.9400 ;
    END
  END sig[1]
  PIN sig[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 65.1400 157.2500 65.2800 ;
    END
  END sig[0]
  PIN speed[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 153.6500 0.5000 153.7900 ;
    END
  END speed[9]
  PIN speed[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 136.5700 0.5000 136.7100 ;
    END
  END speed[8]
  PIN speed[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 119.4900 0.5000 119.6300 ;
    END
  END speed[7]
  PIN speed[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 102.4100 0.5000 102.5500 ;
    END
  END speed[6]
  PIN speed[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 85.3300 0.5000 85.4700 ;
    END
  END speed[5]
  PIN speed[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 68.2500 0.5000 68.3900 ;
    END
  END speed[4]
  PIN speed[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 51.1700 0.5000 51.3100 ;
    END
  END speed[3]
  PIN speed[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 34.0900 0.5000 34.2300 ;
    END
  END speed[2]
  PIN speed[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 17.0100 0.5000 17.1500 ;
    END
  END speed[1]
  PIN speed[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 -0.0700 0.5000 0.0700 ;
    END
  END speed[0]
  PIN TCK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 125.6950 157.2500 125.8350 ;
    END
  END TCK
  PIN scan_done
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 130.3550 157.2500 130.4950 ;
    END
  END scan_done
  PIN over
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 135.0100 157.2500 135.1500 ;
    END
  END over
  PIN test_se
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 139.6700 157.2500 139.8100 ;
    END
  END test_se
  PIN digi_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 144.3300 157.2500 144.4700 ;
    END
  END digi_out
  PIN sub_rst
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 148.9850 157.2500 149.1250 ;
    END
  END sub_rst
  PIN base_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 156.7500 153.6450 157.2500 153.7850 ;
    END
  END base_clk
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER M5 ;
        RECT 154.2500 142.6000 157.2500 145.6000 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 142.6000 3.0000 145.6000 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.2500 8.1200 157.2500 11.1200 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 8.1200 3.0000 11.1200 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.9600 150.7200 148.9600 153.7200 ;
    END
    PORT
      LAYER M4 ;
        RECT 145.9600 0.0000 148.9600 3.0000 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.1200 150.7200 11.1200 153.7200 ;
    END
    PORT
      LAYER M4 ;
        RECT 8.1200 0.0000 11.1200 3.0000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER M5 ;
        RECT 154.2500 147.6000 157.2500 150.6000 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 147.6000 3.0000 150.6000 ;
    END
    PORT
      LAYER M5 ;
        RECT 154.2500 3.1200 157.2500 6.1200 ;
    END
    PORT
      LAYER M5 ;
        RECT 0.0000 3.1200 3.0000 6.1200 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.9600 150.7200 153.9600 153.7200 ;
    END
    PORT
      LAYER M4 ;
        RECT 150.9600 0.0000 153.9600 3.0000 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.1200 150.7200 6.1200 153.7200 ;
    END
    PORT
      LAYER M4 ;
        RECT 3.1200 0.0000 6.1200 3.0000 ;
    END
  END VSS
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 157.2500 153.7200 ;
    LAYER M2 ;
      RECT 147.5850 151.7200 155.6800 153.7200 ;
      RECT 136.3550 151.7200 144.4450 153.7200 ;
      RECT 125.1200 151.7200 133.2150 153.7200 ;
      RECT 113.8900 151.7200 121.9800 153.7200 ;
      RECT 102.6600 151.7200 110.7500 153.7200 ;
      RECT 91.4250 151.7200 99.5200 153.7200 ;
      RECT 80.1950 151.7200 88.2850 153.7200 ;
      RECT 68.9600 151.7200 77.0550 153.7200 ;
      RECT 57.7300 151.7200 65.8200 153.7200 ;
      RECT 46.5000 151.7200 54.5900 153.7200 ;
      RECT 35.2650 151.7200 43.3600 153.7200 ;
      RECT 24.0350 151.7200 32.1250 153.7200 ;
      RECT 12.8000 151.7200 20.8950 153.7200 ;
      RECT 1.5700 151.7200 9.6600 153.7200 ;
      RECT 0.0000 2.0000 157.2500 151.7200 ;
      RECT 150.5400 0.0000 155.6750 2.0000 ;
      RECT 142.2600 0.0000 147.4000 2.0000 ;
      RECT 133.9850 0.0000 139.1200 2.0000 ;
      RECT 125.7100 0.0000 130.8450 2.0000 ;
      RECT 117.4350 0.0000 122.5700 2.0000 ;
      RECT 109.1600 0.0000 114.2950 2.0000 ;
      RECT 100.8800 0.0000 106.0200 2.0000 ;
      RECT 92.6050 0.0000 97.7400 2.0000 ;
      RECT 84.3300 0.0000 89.4650 2.0000 ;
      RECT 76.0550 0.0000 81.1900 2.0000 ;
      RECT 67.7800 0.0000 72.9150 2.0000 ;
      RECT 59.5000 0.0000 64.6400 2.0000 ;
      RECT 51.2250 0.0000 56.3600 2.0000 ;
      RECT 42.9500 0.0000 48.0850 2.0000 ;
      RECT 34.6750 0.0000 39.8100 2.0000 ;
      RECT 26.4000 0.0000 31.5350 2.0000 ;
      RECT 18.1200 0.0000 23.2600 2.0000 ;
      RECT 9.8450 0.0000 14.9800 2.0000 ;
      RECT 1.5700 0.0000 6.7050 2.0000 ;
    LAYER M3 ;
      RECT 2.0000 152.1500 155.2500 153.7200 ;
      RECT 0.0000 152.1450 155.2500 152.1500 ;
      RECT 0.0000 150.6250 157.2500 152.1450 ;
      RECT 0.0000 147.4850 155.2500 150.6250 ;
      RECT 0.0000 145.9700 157.2500 147.4850 ;
      RECT 0.0000 142.8300 155.2500 145.9700 ;
      RECT 0.0000 141.3100 157.2500 142.8300 ;
      RECT 0.0000 138.2100 155.2500 141.3100 ;
      RECT 2.0000 138.1700 155.2500 138.2100 ;
      RECT 2.0000 136.6500 157.2500 138.1700 ;
      RECT 2.0000 135.0700 155.2500 136.6500 ;
      RECT 0.0000 133.5100 155.2500 135.0700 ;
      RECT 0.0000 131.9950 157.2500 133.5100 ;
      RECT 0.0000 128.8550 155.2500 131.9950 ;
      RECT 0.0000 127.3350 157.2500 128.8550 ;
      RECT 0.0000 124.1950 155.2500 127.3350 ;
      RECT 0.0000 122.6800 157.2500 124.1950 ;
      RECT 0.0000 121.1300 155.2500 122.6800 ;
      RECT 2.0000 119.5400 155.2500 121.1300 ;
      RECT 2.0000 118.0200 157.2500 119.5400 ;
      RECT 2.0000 117.9900 155.2500 118.0200 ;
      RECT 0.0000 114.8800 155.2500 117.9900 ;
      RECT 0.0000 113.3600 157.2500 114.8800 ;
      RECT 0.0000 110.2200 155.2500 113.3600 ;
      RECT 0.0000 108.7050 157.2500 110.2200 ;
      RECT 0.0000 105.5650 155.2500 108.7050 ;
      RECT 0.0000 104.0500 157.2500 105.5650 ;
      RECT 2.0000 104.0450 157.2500 104.0500 ;
      RECT 2.0000 100.9100 155.2500 104.0450 ;
      RECT 0.0000 100.9050 155.2500 100.9100 ;
      RECT 0.0000 99.3900 157.2500 100.9050 ;
      RECT 0.0000 96.2500 155.2500 99.3900 ;
      RECT 0.0000 94.7300 157.2500 96.2500 ;
      RECT 0.0000 91.5900 155.2500 94.7300 ;
      RECT 0.0000 90.0700 157.2500 91.5900 ;
      RECT 0.0000 86.9700 155.2500 90.0700 ;
      RECT 2.0000 86.9300 155.2500 86.9700 ;
      RECT 2.0000 85.4150 157.2500 86.9300 ;
      RECT 2.0000 83.8300 155.2500 85.4150 ;
      RECT 0.0000 82.2750 155.2500 83.8300 ;
      RECT 0.0000 80.7550 157.2500 82.2750 ;
      RECT 0.0000 77.6150 155.2500 80.7550 ;
      RECT 0.0000 76.1000 157.2500 77.6150 ;
      RECT 0.0000 72.9600 155.2500 76.1000 ;
      RECT 0.0000 71.4400 157.2500 72.9600 ;
      RECT 0.0000 69.8900 155.2500 71.4400 ;
      RECT 2.0000 68.3000 155.2500 69.8900 ;
      RECT 2.0000 66.7800 157.2500 68.3000 ;
      RECT 2.0000 66.7500 155.2500 66.7800 ;
      RECT 0.0000 63.6400 155.2500 66.7500 ;
      RECT 0.0000 62.1250 157.2500 63.6400 ;
      RECT 0.0000 58.9850 155.2500 62.1250 ;
      RECT 0.0000 57.4650 157.2500 58.9850 ;
      RECT 0.0000 54.3250 155.2500 57.4650 ;
      RECT 0.0000 52.8100 157.2500 54.3250 ;
      RECT 2.0000 49.6700 155.2500 52.8100 ;
      RECT 0.0000 48.1500 157.2500 49.6700 ;
      RECT 0.0000 45.0100 155.2500 48.1500 ;
      RECT 0.0000 43.4900 157.2500 45.0100 ;
      RECT 0.0000 40.3500 155.2500 43.4900 ;
      RECT 0.0000 38.8350 157.2500 40.3500 ;
      RECT 0.0000 35.7300 155.2500 38.8350 ;
      RECT 2.0000 35.6950 155.2500 35.7300 ;
      RECT 2.0000 34.1750 157.2500 35.6950 ;
      RECT 2.0000 32.5900 155.2500 34.1750 ;
      RECT 0.0000 31.0350 155.2500 32.5900 ;
      RECT 0.0000 29.5200 157.2500 31.0350 ;
      RECT 0.0000 26.3800 155.2500 29.5200 ;
      RECT 0.0000 24.8600 157.2500 26.3800 ;
      RECT 0.0000 21.7200 155.2500 24.8600 ;
      RECT 0.0000 20.2000 157.2500 21.7200 ;
      RECT 0.0000 18.6500 155.2500 20.2000 ;
      RECT 2.0000 17.0600 155.2500 18.6500 ;
      RECT 2.0000 15.5450 157.2500 17.0600 ;
      RECT 2.0000 15.5100 155.2500 15.5450 ;
      RECT 0.0000 12.4050 155.2500 15.5100 ;
      RECT 0.0000 10.8850 157.2500 12.4050 ;
      RECT 0.0000 7.7450 155.2500 10.8850 ;
      RECT 0.0000 6.2300 157.2500 7.7450 ;
      RECT 0.0000 3.0900 155.2500 6.2300 ;
      RECT 0.0000 1.5700 157.2500 3.0900 ;
      RECT 2.0000 0.0000 155.2500 1.5700 ;
    LAYER M4 ;
      RECT 155.4600 149.2200 157.2500 153.7200 ;
      RECT 12.6200 149.2200 144.4600 153.7200 ;
      RECT 0.0000 149.2200 1.6200 153.7200 ;
      RECT 0.0000 4.5000 157.2500 149.2200 ;
      RECT 155.4600 0.0000 157.2500 4.5000 ;
      RECT 12.6200 0.0000 144.4600 4.5000 ;
      RECT 0.0000 0.0000 1.6200 4.5000 ;
    LAYER M5 ;
      RECT 0.0000 152.1000 157.2500 153.7200 ;
      RECT 4.5000 141.1000 152.7500 152.1000 ;
      RECT 0.0000 12.6200 157.2500 141.1000 ;
      RECT 4.5000 1.6200 152.7500 12.6200 ;
      RECT 0.0000 0.0000 157.2500 1.6200 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 157.2500 153.7200 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 157.2500 153.7200 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 157.2500 153.7200 ;
    LAYER M9 ;
      RECT 0.0000 0.0000 157.2500 153.7200 ;
  END
END BISG_TOP

END LIBRARY
